/*
*   Copyright 2016 Purdue University
*
*   Licensed under the Apache License, Version 2.0 (the "License");
*   you may not use this file except in compliance with the License.
*   You may obtain a copy of the License at
*
*       http://www.apache.org/licenses/LICENSE-2.0
*
*   Unless required by applicable law or agreed to in writing, software
*   distributed under the License is distributed on an "AS IS" BASIS,
*   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
*   See the License for the specific language governing permissions and
*   limitations under the License.
*
*
*   Filename:     cpu_tracker.sv
*
*   Created by:   Jacob R. Stevens
*   Email:        steven69@purdue.edu
*   Date Created: 06/27/2016
*   Description:  Prints out a trace of the cpu executing that can be
*                 compared against the trace generated by the ISS

    Updated by:   Anusyua Nallathambi, Ansh Patel
    Date: 09/06/2024
*/

`define TRACE_FILE_NAME "cpu_trace.log"

`include "cpu_types_pkg.vh"
import cpu_types_pkg::*;

module cpu_tracker_rv32(
  input logic CLK,
  input logic wb_stall,
  input logic dhit,
  input logic[FUNC3_W-1:0] funct_3,
  input logic[FUNC7_W-1:0] funct_7,
  input opcode_t opcode,
  input regbits_t rs1,
  input regbits_t rs2,
  input regbits_t wsel,
  input word_t instr,
  input word_t pc,
  input word_t next_pc_val,
  input word_t branch_addr,
  input word_t jump_addr,
  input word_t imm,
  input logic [19:0] lui_pre_shift,
  input word_t store_dat,
  input word_t reg_dat,
  input word_t load_dat,
  input word_t dat_addr
);

  parameter CPUID = 0;

  integer fptr, halt_written;
  string instr_mnemonic, output_str, operands, temp_str, halt_temp_str;
  string rs1_str, rs2_str, ram_str, lw_str, halt_output_str, dest_str;
  opcode_t last_opcode;
  funct3_r_t funct3_r;
  funct3_i_t funct3_i;
  funct3_ld_i_t funct3_ld_i;
  funct3_s_t funct3_s;
  funct7_r_t funct7_r;
  funct7_srla_r_t funct7_srla_r;
  funct3_b_t funct3_b;
  funct5_atomic_t funct5;

  initial begin: INIT_FILE
    fptr = $fopen(`TRACE_FILE_NAME, "w");
    halt_written = 0;
  end

  always_comb begin
    rs1_str    = registerAssign(rs1);
    rs2_str    = registerAssign(rs2);
    dest_str  = registerAssign(wsel);
  end

  always_comb begin
    case (opcode)
      RTYPE: $sformat(operands, "%s, %s, %s", dest_str, rs1_str, rs2_str);
      ITYPE: 
      begin
        case(funct3_i_t'(funct_3))
          SRLI_SRAI, SLLI: $sformat(operands, "%s, %s, %d", dest_str, rs1_str, (imm[4:0]));
          default: $sformat(operands, "%s, %s, %d", dest_str, rs1_str, signed'(imm));
        endcase
      end
      LR_SC,ITYPE_LW: $sformat(operands, "%s, %d(%s)", dest_str, signed'(imm), rs1_str);
      STYPE: $sformat(operands, "%s, %d(%s)", rs2_str, signed'(imm), rs1_str);
      JALR: $sformat(operands, "%s, %s, %d", dest_str, rs1_str, signed'(imm));
      BTYPE: $sformat(operands, "%s, %s, %X", rs1_str, rs2_str, branch_addr);
      JAL: $sformat(operands, "%s, %X", dest_str, jump_addr);
      LUI:   $sformat(operands,"%s, %d", dest_str, lui_pre_shift);
      AUIPC: $sformat(operands,"%s, %d", dest_str, lui_pre_shift);
      HALT:  $sformat(operands, "");
    endcase
  end

  always_comb begin
    case (opcode)
      JAL:      instr_mnemonic = "JAL";
      JALR:      instr_mnemonic = "JALR";
      BTYPE:
      begin
        case(funct3_b_t'(funct_3))
          BEQ:      instr_mnemonic = "BEQ";
          BNE:      instr_mnemonic = "BNE";
          BLT:      instr_mnemonic = "BLT";
          BGE:      instr_mnemonic = "BGE";
          BLTU:     instr_mnemonic = "BLTU";
          BGEU:     instr_mnemonic = "BGEU";
        endcase
      end
      STYPE:
      begin
        case(funct3_s_t'(funct_3))
          SB:       instr_mnemonic = "SB";
          SH:       instr_mnemonic = "SH";
          SW:       instr_mnemonic = "SW";
        endcase
      end
      ITYPE_LW:
      begin
        case(funct3_ld_i_t'(funct_3))
          LB:       instr_mnemonic = "LB";
          LH:       instr_mnemonic = "LH";
          LW:       instr_mnemonic = "LW";
          LBU:      instr_mnemonic = "LBU";
          LHU:      instr_mnemonic = "LHU";
        endcase
      end
      LR_SC:
      begin
        case(funct5_atomic_t'(funct_7[4:0]))
          LR:       instr_mnemonic = "LR.W";
          SC:       instr_mnemonic = "SC.W";
        endcase
      end
      ITYPE:
      begin
        case(funct3_i_t'(funct_3))
          ADDI:     instr_mnemonic = "ADDI";
          SLTI:     instr_mnemonic = "SLTI";
          SLTIU:    instr_mnemonic = "SLTIU";
          ANDI:     instr_mnemonic = "ANDI";
          ORI:      instr_mnemonic = "ORI";
          XORI:     instr_mnemonic = "XORI";
          SLLI:     instr_mnemonic = "SLLI";
          SRLI_SRAI:    
          begin
            case(funct7_srla_r_t'(funct_7))
              SRA: instr_mnemonic = "SRAI";
              SRL: instr_mnemonic = "SRLI";
            endcase
          end
        endcase
      end
      LUI:      instr_mnemonic = "LUI";
      AUIPC:   instr_mnemonic = "AUIPC";
      HALT:     instr_mnemonic = "HALT";
      RTYPE: begin
        case(funct3_r_t'(funct_3))
          SLL:  instr_mnemonic = "SLL";
          SRL_SRA:
          begin
            case(funct7_srla_r_t'(funct_7))
              SRA: instr_mnemonic = "SRA";
              SRL: instr_mnemonic = "SRL";
            endcase
          end
          ADD:  instr_mnemonic = "ADD";
          SUB:  instr_mnemonic = "SUB";
          AND:  instr_mnemonic = "AND";
          OR:   instr_mnemonic = "OR";
          XOR:  instr_mnemonic = "XOR";
          SLT:  instr_mnemonic = "SLT";
          SLTU: instr_mnemonic = "SLTU";
        endcase
      end
      default:  instr_mnemonic = "xxx";
    endcase
  end

  function string registerAssign(input logic [4:0] register);
    case (register)
      5'd0:   registerAssign = "R0";
      5'd1:   registerAssign = "R1";
      5'd2:   registerAssign = "R2";
      5'd3:   registerAssign = "R3";
      5'd4:   registerAssign = "R4";
      5'd5:   registerAssign = "R5";
      5'd6:   registerAssign = "R6";
      5'd7:   registerAssign = "R7";
      5'd8:   registerAssign = "R8";
      5'd9:   registerAssign = "R9";
      5'd10:  registerAssign = "R10";
      5'd11:  registerAssign = "R11";
      5'd12:  registerAssign = "R12";
      5'd13:  registerAssign = "R13";
      5'd14:  registerAssign = "R14";
      5'd15:  registerAssign = "R15";
      5'd16:  registerAssign = "R16";
      5'd17:  registerAssign = "R17";
      5'd18:  registerAssign = "R18";
      5'd19:  registerAssign = "R19";
      5'd20:  registerAssign = "R20";
      5'd21:  registerAssign = "R21";
      5'd22:  registerAssign = "R22";
      5'd23:  registerAssign = "R23";
      5'd24:  registerAssign = "R24";
      5'd25:  registerAssign = "R25";
      5'd26:  registerAssign = "R26";
      5'd27:  registerAssign = "R27";
      5'd28:  registerAssign = "R28";
      5'd29:  registerAssign = "R29";
      5'd30:  registerAssign = "R30";
      5'd31:  registerAssign = "R31";
    endcase
  endfunction

  always_ff @ (posedge CLK) begin
    if (dhit) begin
        if (last_opcode == ITYPE_LW) begin
          $sformat(temp_str, "%X (Core %d): %X", pc, CPUID + 1, instr);
          $sformat(temp_str, "%s %s %s\n", temp_str, instr_mnemonic, operands);
          $sformat(ram_str, "    [word read");
          $sformat(ram_str, "%s from %x]\n", ram_str, {16'h0, dat_addr[15:0]});
          $sformat(ram_str, "%s    %s", ram_str, dest_str);
          $sformat(ram_str, "%s <-- %x\n", ram_str, load_dat);
          $sformat(lw_str, "%s%s\n", temp_str, ram_str);
          $fwrite(fptr, lw_str);
        end
    end
  end

  always_ff @ (posedge CLK) begin
    if (!wb_stall)
      last_opcode <= opcode;
  end

  always_ff @ (posedge CLK) begin
    if (!wb_stall && instr != 0) begin
      $sformat(temp_str, "%X (Core %d): %X", pc, CPUID + 1, instr);
      $sformat(temp_str, "%s %s %s\n", temp_str, instr_mnemonic, operands);
      $sformat(temp_str, "%s    PC <-- %X\n", temp_str, next_pc_val);
      case(opcode)
        RTYPE: 
        begin
          case(funct3_r_t'(funct_3))
            SLL:  $sformat(temp_str, "%s    %s <-- %x\n", temp_str, dest_str, reg_dat);
            SRL_SRA:
            begin
              case(funct7_srla_r_t'(funct_7))
                SRA: $sformat(temp_str, "%s    %s <-- %x\n", temp_str, dest_str, reg_dat);
                SRL: $sformat(temp_str, "%s    %s <-- %x\n", temp_str, dest_str, reg_dat);
              endcase
            end
            ADD, SUB, AND, OR, XOR, SLT, SLTU: $sformat(temp_str, "%s    %s <-- %x\n", temp_str, dest_str, reg_dat);
          endcase
        end
        ITYPE:
        begin
          case(funct3_i_t'(funct_3))
            default: $sformat(temp_str, "%s    %s <-- %x\n", temp_str, dest_str, reg_dat);
          endcase
        end
        BTYPE:
        begin
          case(funct3_b_t'(funct_3))
            default: $sformat(temp_str, "%s    %s <-- %x\n", temp_str, dest_str, reg_dat);
          endcase
        end
        JAL, JALR: $sformat(temp_str, "%s    %s <-- %x\n", temp_str, dest_str, reg_dat);
        LUI:  $sformat(temp_str, "%s    %s <-- %x\n", temp_str, dest_str, {lui_pre_shift, 12'b0});
        AUIPC:  $sformat(temp_str, "%s    %s <-- %x\n", temp_str, dest_str, pc+(lui_pre_shift<<12));
        STYPE: begin
              $sformat(temp_str,"%s    [%x]",temp_str,{16'h0, dat_addr[15:0]});
              $sformat(temp_str, "%s <-- %x\n", temp_str, store_dat);
        end
        //TODO: add atomic instructions
        default: $sformat(temp_str, "");
      endcase
      $sformat(output_str, "%s\n", temp_str);
      $fwrite(fptr, output_str);
    end
  end

  final begin: CLOSE_FILE
    $fclose(fptr);
  end

endmodule
